module lab7_tb();
  reg clk,reset;


lab7_top DUT(clk,reset);
initial begin 
	clk = 0;
	reset = 1;
	#5;
	clk = 1;
	#5;
	clk = 0;
	#5;
	reset = 0; 
	clk = 1;
	#5;
	clk = 0; 
	#5;
	clk = 1;
	#5;
	clk = 0; 
	#5;
	clk = 1;
	#5;
	clk = 0; 
	#5;
	clk = 1;
	#5;
	clk = 0; 
         #5;
	clk = 1;
	#5;
	clk = 0; 
	#5;
	clk = 1;
	#5;
clk = 0; 
	#5;
	clk = 1;
	#5;
	
clk = 0; 
	#5;
	clk = 1;
	#5;
	
clk = 0; 
	#5;
	clk = 1;
	#5;
	
clk = 0; 
	#5;
	clk = 1;
	#5;
clk = 0; 
	#5;
	clk = 1;
	#5;
	
clk = 0; 
	#5;
	clk = 1;
	#5;
	
clk = 0; 
	#5;
	clk = 1;
	#5;
	
	
clk = 0; 
	#5;
	clk = 1;
	#5;
	
clk = 0; 
	#5;
	clk = 1;
	#5;
	
clk = 0; 
	#5;
	clk = 1;
	#5;
	
	clk = 0; 
	#5;
	clk = 1;
	#5;
	
clk = 0; 
	#5;
	clk = 1;
	#5;
	
clk = 0; 
	#5;
	clk = 1;
	#5;
	
	clk = 0; 
	#5;
	clk = 1;
	#5;
	
clk = 0; 
	#5;
	clk = 1;
	#5;
	
clk = 0; 
	#5;
	clk = 1;
	#5;
	
	clk = 0; 
	#5;
	clk = 1;
	#5;
	
clk = 0; 
	#5;
	clk = 1;
	#5;
	
clk = 0; 
	#5;
	clk = 1;
	#5;
	
clk = 0; 
	#5;
	clk = 1;
	#5;
	
clk = 0; 
	#5;
	clk = 1;
	#5;
	
clk = 0; 
	#5;
	clk = 1;
	#5;
	
	
clk = 0; 
	#5;
	clk = 1;
	#5;
	
clk = 0; 
	#5;
	clk = 1;
	#5;
	
clk = 0; 
	#5;
	clk = 1;
	#5;
	
	clk = 0; 
	#5;
	clk = 1;
	#5;
	clk = 0; 
	#5;
	clk = 1;
	#5;
	
	clk = 0; 
	#5;
	clk = 1;
	#5;
clk = 0; 
	#5;
	clk = 1;
	#5;
	clk = 0; 
	#5;
	clk = 1;
	#5;
	
	clk = 0; 
	#5;
	clk = 1;
	#5;
clk = 0; 
	#5;
	clk = 1;
	#5;
	clk = 0; 
	#5;
	clk = 1;
	#5;
	
	clk = 0; 
	#5;
	clk = 1;
	#5;
clk = 0; 
	#5;
	clk = 1;
	#5;
	clk = 0; 
	#5;
	clk = 1;
	#5;
	
	clk = 0; 
	#5;
	clk = 1;
	#5;
clk = 0; 
	#5;
	clk = 1;
	#5;
	clk = 0; 
	#5;
	clk = 1;
	#5;
	
	clk = 0; 
	#5;
	clk = 1;
	#5;
clk = 0; 
	#5;
	clk = 1;
	#5;
	clk = 0; 
	#5;
	clk = 1;
	#5;
	
	clk = 0; 
	#5;
	clk = 1;
	#5;
clk = 0; 
	#5;
	clk = 1;
	#5;
	clk = 0; 
	#5;
	clk = 1;
	#5;
	
	clk = 0; 
	#5;
	clk = 1;
	#5;
clk = 0; 
	#5;
	clk = 1;
	#5;
	clk = 0; 
	#5;
	clk = 1;
	#5;
	
	clk = 0; 
	#5;
	clk = 1;
	#5;
clk = 0; 
	#5;
	clk = 1;
	#5;
	clk = 0; 
	#5;
	clk = 1;
	#5;
	
	clk = 0; 
	#5;
	clk = 1;
	#5;
clk = 0; 
	#5;
	clk = 1;
	#5;
	clk = 0; 
	#5;
	clk = 1;
	#5;
	
	clk = 0; 
	#5;
	clk = 1;
	#5;
clk = 0; 
	#5;
	clk = 1;
	#5;
	clk = 0; 
	#5;
	clk = 1;
	#5;
	
	clk = 0; 
	#5;
	clk = 1;
	#5;
clk = 0; 
	#5;
	clk = 1;
	#5;
	clk = 0; 
	#5;
	clk = 1;
	#5;
	
	clk = 0; 
	#5;
	clk = 1;
	#5;
clk = 0; 
	#5;
	clk = 1;
	#5;
	clk = 0; 
	#5;
	clk = 1;
	#5;
	
	clk = 0; 
	#5;
	clk = 1;
	#5;
	clk = 0; 
	#5;
	clk = 1;
	#5;
	
	clk = 0; 
	#5;
	clk = 1;
	#5;
	clk = 0; 
	#5;
	clk = 1;
	#5;
	clk = 0; 
	#5;
	clk = 1;
	#5;
	
	clk = 0; 
	#5;
	clk = 1;
	#5;
	clk = 0; 
	#5;
	clk = 1;
	#5;
	clk = 0; 
	#5;
	clk = 1;
	#5;
	
	clk = 0; 
	#5;
	clk = 1;
	#5;
	clk = 0; 
	#5;
	clk = 1;
	#5;
	clk = 0; 
	#5;
	clk = 1;
	#5;
	
	clk = 0; 
	#5;
	clk = 1;
	#5;
	clk = 0; 
	#5;
	clk = 1;
	#5;
	clk = 0; 
	#5;
	clk = 1;
	#5;
	
	clk = 0; 
	#5;
	clk = 1;
	#5;


	clk = 0; 
	#5;
	clk = 1;
	#5;
	clk = 0; 
	#5;
	clk = 1;
	#5;
	
	clk = 0; 
	#5;
	clk = 1;
	#5;

	$stop;

end 


endmodule
